    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   LoadSavePref+Position   xyz      �f�  �@@%�>